--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Alutosel is
    Port ( ALU : in  STD_LOGIC_VECTOR (4 downto 0);
           sel : out  STD_LOGIC_VECTOR (1 downto 0));
end Alutosel;

architecture Behavioral of Alutosel is

begin


end Behavioral;

